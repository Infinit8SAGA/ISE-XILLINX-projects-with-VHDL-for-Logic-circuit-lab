----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    21:13:37 05/08/2025 
-- Design Name: 
-- Module Name:    main - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


entity main is
	port (
		T : in STD_LOGIC; -- ????? ????
		CLK : in STD_LOGIC;-- ?????? ????
		RESET : in STD_LOGIC;--????? ????
		Q : out STD_LOGIC-- ????? ???? ????
	);
end main;

architecture Behavioral of main is
	signal internal_state : STD_LOGIC := '0'; -- ???? ????? ??????? ????? ???
begin
	process(CLK, RESET)--???? ???? ?? ???? ? ????
	begin
		if RESET = '1' then -- ??? ???? ?????? ??????
			internal_state <= '0';-- ???? ??????
		elsif rising_edge(CLK) then-- ??? ????????? ????
			if T = '1' then --???? ?? ???? ????
				internal_state <= not internal_state;--????? ????
			end if;	--??? ?? ????? ??? ???? ???? ??? ?????
		end if;	
	end process;
	Q <= internal_state;-- ?????? ?????
end Behavioral;

